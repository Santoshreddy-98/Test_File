VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;


MANUFACTURINGGRID 0.005 ;

MACRO BUFFSGD3BWP30P140HVT
    CLASS CORE ;
    FOREIGN BUFFSGD3BWP30P140HVT 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 0.900 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120900 ;
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.145 0.675 0.755 ;
        RECT  0.605 0.145 0.625 0.340 ;
        RECT  0.605 0.545 0.625 0.755 ;
        RECT  0.375 0.290 0.605 0.340 ;
        RECT  0.375 0.545 0.605 0.595 ;
        RECT  0.325 0.145 0.375 0.340 ;
        RECT  0.325 0.545 0.375 0.745 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.385 0.170 0.480 ;
        RECT  0.035 0.345 0.105 0.555 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 -0.075 0.700 0.075 ;
        RECT  0.450 -0.075 0.530 0.240 ;
        RECT  0.250 -0.075 0.450 0.075 ;
        RECT  0.170 -0.075 0.250 0.170 ;
        RECT  0.000 -0.075 0.170 0.075 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.825 0.700 0.975 ;
        RECT  0.455 0.645 0.525 0.975 ;
        RECT  0.250 0.825 0.455 0.975 ;
        RECT  0.170 0.735 0.250 0.975 ;
        RECT  0.000 0.825 0.170 0.975 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT  0.610 0.170 0.650 0.210 ;
        RECT  0.610 0.280 0.650 0.320 ;
        RECT  0.610 0.580 0.650 0.620 ;
        RECT  0.610 0.690 0.650 0.730 ;
        RECT  0.535 0.410 0.575 0.450 ;
        RECT  0.470 0.085 0.510 0.125 ;
        RECT  0.470 0.195 0.510 0.235 ;
        RECT  0.470 0.660 0.510 0.700 ;
        RECT  0.470 0.770 0.510 0.810 ;
        RECT  0.400 0.405 0.440 0.445 ;
        RECT  0.330 0.165 0.370 0.205 ;
        RECT  0.330 0.275 0.370 0.315 ;
        RECT  0.330 0.575 0.370 0.615 ;
        RECT  0.330 0.685 0.370 0.725 ;
        RECT  0.260 0.405 0.300 0.445 ;
        RECT  0.190 0.120 0.230 0.160 ;
        RECT  0.190 0.745 0.230 0.785 ;
        RECT  0.120 0.410 0.160 0.450 ;
        RECT  0.050 0.195 0.090 0.235 ;
        RECT  0.050 0.665 0.090 0.705 ;
        LAYER M1 ;
        RECT  0.505 0.390 0.575 0.480 ;
        RECT  0.275 0.390 0.505 0.450 ;
        RECT  0.225 0.230 0.275 0.685 ;
        RECT  0.105 0.230 0.225 0.280 ;
        RECT  0.105 0.635 0.225 0.685 ;
        RECT  0.035 0.180 0.105 0.280 ;
        RECT  0.035 0.635 0.105 0.735 ;
    END
END BUFFSGD3BWP30P140HVT

MACRO SDFQOPPSBSGD1BWP30P140HVT
    CLASS CORE ;
    FOREIGN SDFQOPPSBSGD1BWP30P140HVT 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 0.900 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.006000 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M2 ;
        RECT  0.595 0.375 0.905 0.425 ;
        VIA  0.685 0.4 VIA12_square ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.018450 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.785 0.255 0.835 0.625 ;
        RECT  0.600 0.255 0.785 0.305 ;
        RECT  0.465 0.575 0.785 0.625 ;
        RECT  0.520 0.255 0.600 0.325 ;
        RECT  0.385 0.475 0.465 0.625 ;
        RECT  0.175 0.575 0.385 0.625 ;
        RECT  0.125 0.445 0.175 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.052700 ;
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  3.145 0.125 3.195 0.755 ;
        RECT  3.125 0.125 3.145 0.335 ;
        RECT  3.125 0.545 3.145 0.755 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.012450 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.225 0.375 0.335 0.525 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.012000 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M2 ;
        RECT  0.830 0.475 1.140 0.525 ;
        VIA  0.945 0.5 VIA12_square ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.050 -0.075 3.220 0.075 ;
        RECT  2.970 -0.075 3.050 0.235 ;
        RECT  2.760 -0.075 2.970 0.075 ;
        RECT  2.710 -0.075 2.760 0.175 ;
        RECT  2.195 -0.075 2.710 0.075 ;
        RECT  2.145 -0.075 2.195 0.175 ;
        RECT  1.925 -0.075 2.145 0.075 ;
        RECT  1.855 -0.075 1.925 0.160 ;
        RECT  1.075 -0.075 1.855 0.075 ;
        RECT  1.025 -0.075 1.075 0.175 ;
        RECT  0.795 -0.075 1.025 0.075 ;
        RECT  0.745 -0.075 0.795 0.175 ;
        RECT  0.250 -0.075 0.745 0.075 ;
        RECT  0.170 -0.075 0.250 0.125 ;
        RECT  0.000 -0.075 0.170 0.075 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.035 0.825 3.220 0.975 ;
        RECT  2.985 0.635 3.035 0.975 ;
        RECT  2.760 0.825 2.985 0.975 ;
        RECT  2.710 0.730 2.760 0.975 ;
        RECT  2.195 0.825 2.710 0.975 ;
        RECT  2.145 0.685 2.195 0.975 ;
        RECT  1.930 0.825 2.145 0.975 ;
        RECT  1.850 0.780 1.930 0.975 ;
        RECT  1.075 0.825 1.850 0.975 ;
        RECT  1.025 0.725 1.075 0.975 ;
        RECT  0.795 0.825 1.025 0.975 ;
        RECT  0.745 0.725 0.795 0.975 ;
        RECT  0.230 0.825 0.745 0.975 ;
        RECT  0.180 0.720 0.230 0.975 ;
        RECT  0.000 0.825 0.180 0.975 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT  3.130 0.155 3.170 0.195 ;
        RECT  3.130 0.265 3.170 0.305 ;
        RECT  3.130 0.570 3.170 0.610 ;
        RECT  3.130 0.680 3.170 0.720 ;
        RECT  3.055 0.400 3.095 0.440 ;
        RECT  2.990 0.080 3.030 0.120 ;
        RECT  2.990 0.190 3.030 0.230 ;
        RECT  2.990 0.665 3.030 0.705 ;
        RECT  2.990 0.775 3.030 0.815 ;
        RECT  2.920 0.405 2.960 0.445 ;
        RECT  2.850 0.125 2.890 0.165 ;
        RECT  2.850 0.735 2.890 0.775 ;
        RECT  2.710 0.105 2.750 0.145 ;
        RECT  2.710 0.755 2.750 0.795 ;
        RECT  2.640 0.480 2.680 0.520 ;
        RECT  2.500 0.385 2.540 0.425 ;
        RECT  2.500 0.555 2.540 0.595 ;
        RECT  2.430 0.130 2.470 0.170 ;
        RECT  2.430 0.715 2.470 0.755 ;
        RECT  2.360 0.300 2.400 0.340 ;
        RECT  2.360 0.545 2.400 0.585 ;
        RECT  2.220 0.560 2.260 0.600 ;
        RECT  2.150 0.105 2.190 0.145 ;
        RECT  2.150 0.720 2.190 0.760 ;
        RECT  2.010 0.125 2.050 0.165 ;
        RECT  2.010 0.735 2.050 0.775 ;
        RECT  1.940 0.560 1.980 0.600 ;
        RECT  1.870 0.105 1.910 0.145 ;
        RECT  1.870 0.780 1.910 0.820 ;
        RECT  1.800 0.265 1.840 0.305 ;
        RECT  1.730 0.125 1.770 0.165 ;
        RECT  1.730 0.725 1.770 0.765 ;
        RECT  1.660 0.460 1.700 0.500 ;
        RECT  1.590 0.125 1.630 0.165 ;
        RECT  1.590 0.735 1.630 0.775 ;
        RECT  1.520 0.360 1.560 0.400 ;
        RECT  1.515 0.575 1.555 0.615 ;
        RECT  1.450 0.140 1.490 0.180 ;
        RECT  1.450 0.735 1.490 0.775 ;
        RECT  1.380 0.405 1.420 0.445 ;
        RECT  1.380 0.575 1.420 0.615 ;
        RECT  1.310 0.125 1.350 0.165 ;
        RECT  1.310 0.735 1.350 0.775 ;
        RECT  1.170 0.280 1.210 0.320 ;
        RECT  1.170 0.560 1.210 0.600 ;
        RECT  1.100 0.410 1.140 0.450 ;
        RECT  1.030 0.105 1.070 0.145 ;
        RECT  1.030 0.755 1.070 0.795 ;
        RECT  0.960 0.410 1.000 0.450 ;
        RECT  0.890 0.155 0.930 0.195 ;
        RECT  0.890 0.265 0.930 0.305 ;
        RECT  0.890 0.595 0.930 0.635 ;
        RECT  0.890 0.705 0.930 0.745 ;
        RECT  0.750 0.105 0.790 0.145 ;
        RECT  0.750 0.755 0.790 0.795 ;
        RECT  0.680 0.445 0.720 0.485 ;
        RECT  0.540 0.280 0.580 0.320 ;
        RECT  0.540 0.445 0.580 0.485 ;
        RECT  0.470 0.145 0.510 0.185 ;
        RECT  0.470 0.715 0.510 0.755 ;
        RECT  0.405 0.475 0.445 0.515 ;
        RECT  0.400 0.285 0.440 0.325 ;
        RECT  0.330 0.145 0.370 0.185 ;
        RECT  0.330 0.705 0.370 0.745 ;
        RECT  0.260 0.400 0.300 0.440 ;
        RECT  0.190 0.085 0.230 0.125 ;
        RECT  0.190 0.755 0.230 0.795 ;
        RECT  0.125 0.475 0.165 0.515 ;
        RECT  0.050 0.125 0.090 0.165 ;
        RECT  0.050 0.735 0.090 0.775 ;
        LAYER M1 ;
        RECT  3.060 0.380 3.095 0.460 ;
        RECT  3.010 0.285 3.060 0.565 ;
        RECT  2.910 0.285 3.010 0.335 ;
        RECT  2.910 0.515 3.010 0.565 ;
        RECT  2.795 0.385 2.960 0.465 ;
        RECT  2.860 0.125 2.910 0.335 ;
        RECT  2.860 0.515 2.910 0.775 ;
        RECT  2.830 0.125 2.860 0.180 ;
        RECT  2.830 0.720 2.860 0.775 ;
        RECT  2.745 0.290 2.795 0.660 ;
        RECT  2.660 0.290 2.745 0.340 ;
        RECT  2.660 0.610 2.745 0.660 ;
        RECT  2.610 0.390 2.695 0.560 ;
        RECT  2.610 0.145 2.660 0.340 ;
        RECT  2.610 0.610 2.660 0.745 ;
        RECT  2.490 0.145 2.610 0.195 ;
        RECT  2.495 0.695 2.610 0.745 ;
        RECT  2.480 0.375 2.560 0.460 ;
        RECT  2.455 0.510 2.560 0.645 ;
        RECT  2.405 0.275 2.505 0.325 ;
        RECT  2.425 0.695 2.495 0.775 ;
        RECT  2.410 0.125 2.490 0.195 ;
        RECT  2.405 0.410 2.480 0.460 ;
        RECT  2.355 0.275 2.405 0.360 ;
        RECT  2.355 0.410 2.405 0.605 ;
        RECT  2.230 0.310 2.355 0.360 ;
        RECT  2.350 0.455 2.355 0.605 ;
        RECT  1.430 0.455 2.350 0.505 ;
        RECT  1.655 0.555 2.280 0.605 ;
        RECT  2.180 0.310 2.230 0.405 ;
        RECT  1.500 0.355 2.180 0.405 ;
        RECT  1.980 0.655 2.095 0.775 ;
        RECT  2.025 0.125 2.070 0.195 ;
        RECT  1.975 0.125 2.025 0.305 ;
        RECT  1.925 0.655 1.980 0.730 ;
        RECT  1.775 0.255 1.975 0.305 ;
        RECT  1.800 0.655 1.855 0.730 ;
        RECT  1.705 0.655 1.800 0.775 ;
        RECT  1.705 0.125 1.790 0.195 ;
        RECT  1.630 0.125 1.705 0.305 ;
        RECT  1.650 0.555 1.655 0.725 ;
        RECT  1.605 0.555 1.650 0.775 ;
        RECT  1.570 0.125 1.630 0.195 ;
        RECT  1.430 0.700 1.605 0.775 ;
        RECT  1.355 0.555 1.555 0.635 ;
        RECT  1.420 0.125 1.520 0.265 ;
        RECT  1.325 0.340 1.430 0.505 ;
        RECT  1.260 0.125 1.370 0.195 ;
        RECT  1.260 0.705 1.370 0.775 ;
        RECT  1.260 0.555 1.355 0.605 ;
        RECT  1.150 0.125 1.260 0.225 ;
        RECT  1.210 0.275 1.260 0.605 ;
        RECT  1.150 0.675 1.260 0.775 ;
        RECT  1.150 0.275 1.210 0.345 ;
        RECT  1.150 0.535 1.210 0.605 ;
        RECT  1.100 0.395 1.160 0.465 ;
        RECT  1.050 0.275 1.100 0.625 ;
        RECT  0.935 0.275 1.050 0.325 ;
        RECT  0.935 0.575 1.050 0.625 ;
        RECT  0.885 0.375 1.000 0.525 ;
        RECT  0.885 0.135 0.935 0.325 ;
        RECT  0.885 0.575 0.935 0.765 ;
        RECT  0.635 0.365 0.735 0.505 ;
        RECT  0.465 0.125 0.685 0.205 ;
        RECT  0.565 0.675 0.675 0.775 ;
        RECT  0.515 0.375 0.585 0.505 ;
        RECT  0.470 0.695 0.565 0.775 ;
        RECT  0.460 0.375 0.515 0.425 ;
        RECT  0.400 0.275 0.460 0.425 ;
        RECT  0.280 0.675 0.420 0.775 ;
        RECT  0.310 0.125 0.405 0.225 ;
        RECT  0.110 0.275 0.400 0.325 ;
        RECT  0.190 0.175 0.310 0.225 ;
        RECT  0.075 0.125 0.110 0.325 ;
        RECT  0.075 0.705 0.110 0.775 ;
        RECT  0.025 0.125 0.075 0.775 ;
        LAYER VIA1 ;
        RECT  3.010 0.475 3.060 0.525 ;
        RECT  2.635 0.475 2.685 0.525 ;
        RECT  2.480 0.575 2.530 0.625 ;
        RECT  2.405 0.275 2.455 0.325 ;
        RECT  2.010 0.675 2.060 0.725 ;
        RECT  1.945 0.255 1.995 0.305 ;
        RECT  1.735 0.675 1.785 0.725 ;
        RECT  1.645 0.230 1.695 0.280 ;
        RECT  1.475 0.700 1.525 0.750 ;
        RECT  1.450 0.175 1.500 0.225 ;
        RECT  1.325 0.375 1.375 0.425 ;
        RECT  1.180 0.175 1.230 0.225 ;
        RECT  1.180 0.675 1.230 0.725 ;
        RECT  1.050 0.375 1.100 0.425 ;
        RECT  0.605 0.145 0.655 0.195 ;
        RECT  0.595 0.685 0.645 0.735 ;
        RECT  0.325 0.175 0.375 0.225 ;
        RECT  0.325 0.675 0.375 0.725 ;
        LAYER M2 ;
        RECT  2.585 0.475 3.110 0.525 ;
        RECT  2.405 0.575 2.580 0.625 ;
        RECT  2.405 0.275 2.505 0.325 ;
        RECT  2.355 0.275 2.405 0.625 ;
        RECT  1.965 0.675 2.110 0.725 ;
        RECT  1.965 0.255 2.035 0.305 ;
        RECT  1.915 0.255 1.965 0.725 ;
        RECT  1.660 0.675 1.835 0.725 ;
        RECT  1.660 0.230 1.740 0.280 ;
        RECT  1.610 0.230 1.660 0.725 ;
        RECT  1.505 0.175 1.555 0.750 ;
        RECT  1.400 0.175 1.505 0.225 ;
        RECT  1.445 0.700 1.505 0.750 ;
        RECT  1.000 0.375 1.425 0.425 ;
        RECT  0.685 0.175 1.260 0.225 ;
        RECT  0.675 0.675 1.260 0.725 ;
        RECT  0.575 0.135 0.685 0.225 ;
        RECT  0.565 0.675 0.675 0.745 ;
        RECT  0.465 0.175 0.515 0.725 ;
        RECT  0.275 0.175 0.465 0.225 ;
        RECT  0.275 0.675 0.465 0.725 ;
    END
END SDFQOPPSBSGD1BWP30P140HVT

MACRO XOR2SGD0BWP30P140
    CLASS CORE ;
    FOREIGN XOR2SGD0BWP30P140 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 0.900 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.026350 ;
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.125 1.095 0.775 ;
        RECT  1.025 0.125 1.045 0.205 ;
        RECT  1.010 0.725 1.045 0.775 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.009300 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M2 ;
        RECT  0.875 0.175 1.035 0.225 ;
        RECT  0.825 0.175 0.875 0.495 ;
        RECT  0.725 0.175 0.825 0.225 ;
        VIA  0.85 0.42 VIA12_square ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M2 ;
        RECT  0.375 0.375 0.445 0.480 ;
        RECT  0.115 0.375 0.375 0.425 ;
        VIA  0.41 0.43 VIA12_square ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.075 1.120 0.075 ;
        RECT  0.875 -0.075 0.945 0.180 ;
        RECT  0.230 -0.075 0.875 0.075 ;
        RECT  0.160 -0.075 0.230 0.180 ;
        RECT  0.000 -0.075 0.160 0.075 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 0.825 1.120 0.975 ;
        RECT  0.885 0.645 0.935 0.975 ;
        RECT  0.235 0.825 0.885 0.975 ;
        RECT  0.185 0.645 0.235 0.975 ;
        RECT  0.000 0.825 0.185 0.975 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT  1.030 0.145 1.070 0.185 ;
        RECT  1.030 0.730 1.070 0.770 ;
        RECT  0.955 0.410 0.995 0.450 ;
        RECT  0.890 0.125 0.930 0.165 ;
        RECT  0.890 0.665 0.930 0.705 ;
        RECT  0.890 0.775 0.930 0.815 ;
        RECT  0.820 0.410 0.860 0.450 ;
        RECT  0.750 0.145 0.790 0.185 ;
        RECT  0.750 0.735 0.790 0.775 ;
        RECT  0.675 0.410 0.715 0.450 ;
        RECT  0.610 0.145 0.650 0.185 ;
        RECT  0.610 0.530 0.650 0.570 ;
        RECT  0.535 0.315 0.575 0.355 ;
        RECT  0.470 0.145 0.510 0.185 ;
        RECT  0.470 0.730 0.510 0.770 ;
        RECT  0.400 0.410 0.440 0.450 ;
        RECT  0.330 0.145 0.370 0.185 ;
        RECT  0.330 0.700 0.370 0.740 ;
        RECT  0.265 0.505 0.305 0.545 ;
        RECT  0.190 0.120 0.230 0.160 ;
        RECT  0.190 0.665 0.230 0.705 ;
        RECT  0.190 0.775 0.230 0.815 ;
        RECT  0.125 0.425 0.165 0.465 ;
        RECT  0.050 0.140 0.090 0.180 ;
        RECT  0.050 0.720 0.090 0.760 ;
        LAYER M1 ;
        RECT  0.925 0.390 0.995 0.575 ;
        RECT  0.875 0.290 0.955 0.340 ;
        RECT  0.565 0.525 0.925 0.575 ;
        RECT  0.825 0.290 0.875 0.475 ;
        RECT  0.805 0.395 0.825 0.475 ;
        RECT  0.730 0.625 0.810 0.775 ;
        RECT  0.775 0.125 0.795 0.205 ;
        RECT  0.665 0.125 0.775 0.355 ;
        RECT  0.175 0.405 0.735 0.455 ;
        RECT  0.495 0.625 0.730 0.675 ;
        RECT  0.605 0.125 0.665 0.205 ;
        RECT  0.105 0.305 0.595 0.355 ;
        RECT  0.445 0.125 0.555 0.255 ;
        RECT  0.375 0.725 0.540 0.775 ;
        RECT  0.445 0.505 0.495 0.675 ;
        RECT  0.245 0.505 0.445 0.555 ;
        RECT  0.280 0.125 0.390 0.255 ;
        RECT  0.325 0.645 0.375 0.775 ;
        RECT  0.125 0.405 0.175 0.485 ;
        RECT  0.075 0.125 0.105 0.355 ;c
        RECT  0.075 0.705 0.105 0.775 ;
        RECT  0.025 0.125 0.075 0.775 ;
        LAYER VIA1 ;
        RECT  0.695 0.305 0.745 0.355 ;
        RECT  0.695 0.625 0.745 0.675 ;
        RECT  0.595 0.525 0.645 0.575 ;
        RECT  0.505 0.175 0.555 0.225 ;
        RECT  0.325 0.675 0.375 0.725 ;
        RECT  0.295 0.175 0.345 0.225 ;
        LAYER M2 ;
        RECT  0.745 0.675 0.800 0.725 ;
        RECT  0.745 0.275 0.765 0.345 ;
        RECT  0.695 0.275 0.745 0.725 ;
        RECT  0.595 0.175 0.645 0.625 ;
        RECT  0.455 0.175 0.595 0.225 ;
        RECT  0.495 0.275 0.545 0.725 ;
        RECT  0.375 0.275 0.495 0.325 ;
        RECT  0.275 0.675 0.495 0.725 ;
        RECT  0.325 0.175 0.375 0.325 ;
        RECT  0.245 0.175 0.325 0.225 ;
    END
END XOR2SGD0BWP30P140


MACRO AN2SGD0BWP30P140
    CLASS CORE ;
    FOREIGN AN2SGD0BWP30P140 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 0.900 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.026350 ;
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.485 0.125 0.535 0.755 ;
        RECT  0.465 0.125 0.485 0.335 ;
        RECT  0.465 0.545 0.485 0.755 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.009300 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.400 0.315 0.470 ;
        RECT  0.230 0.145 0.280 0.470 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.009300 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.245 0.180 0.500 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.395 -0.075 0.560 0.075 ;
        RECT  0.330 -0.075 0.395 0.180 ;
        RECT  0.000 -0.075 0.330 0.075 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.825 0.560 0.975 ;
        RECT  0.310 0.660 0.390 0.975 ;
        RECT  0.110 0.825 0.310 0.975 ;
        RECT  0.030 0.735 0.110 0.975 ;
        RECT  0.000 0.825 0.030 0.975 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT  0.470 0.145 0.510 0.185 ;
        RECT  0.470 0.695 0.510 0.735 ;
        RECT  0.395 0.410 0.435 0.450 ;
        RECT  0.330 0.110 0.370 0.150 ;
        RECT  0.330 0.665 0.370 0.705 ;
        RECT  0.330 0.775 0.370 0.815 ;
        RECT  0.260 0.415 0.300 0.455 ;
        RECT  0.190 0.695 0.230 0.735 ;
        RECT  0.125 0.375 0.165 0.415 ;
        RECT  0.050 0.130 0.090 0.170 ;
        RECT  0.050 0.740 0.090 0.780 ;
        LAYER M1 ;
        RECT  0.415 0.390 0.435 0.470 ;
        RECT  0.365 0.390 0.415 0.610 ;
        RECT  0.245 0.560 0.365 0.610 ;
        RECT  0.205 0.560 0.245 0.755 ;
        RECT  0.185 0.570 0.205 0.755 ;
        RECT  0.075 0.570 0.185 0.620 ;
        RECT  0.075 0.125 0.110 0.175 ;
        RECT  0.025 0.125 0.075 0.620 ;
    END
END AN2SGD0BWP30P140




MACRO OR2SGD1BWP30P140
    CLASS CORE ;
    FOREIGN OR2SGD1BWP30P140 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 0.900 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.052700 ;
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.485 0.125 0.535 0.755 ;
        RECT  0.465 0.125 0.485 0.315 ;
        RECT  0.465 0.555 0.485 0.755 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.014400 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.235 0.345 0.305 0.555 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.014400 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.345 0.155 0.425 ;
        RECT  0.035 0.345 0.105 0.555 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.390 -0.075 0.560 0.075 ;
        RECT  0.310 -0.075 0.390 0.190 ;
        RECT  0.095 -0.075 0.310 0.075 ;
        RECT  0.045 -0.075 0.095 0.175 ;
        RECT  0.000 -0.075 0.045 0.075 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.825 0.560 0.975 ;
        RECT  0.315 0.705 0.385 0.975 ;
        RECT  0.000 0.825 0.315 0.975 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT  0.470 0.145 0.510 0.185 ;
        RECT  0.470 0.255 0.510 0.295 ;
        RECT  0.470 0.575 0.510 0.615 ;
        RECT  0.470 0.685 0.510 0.725 ;
        RECT  0.395 0.400 0.435 0.440 ;
        RECT  0.330 0.145 0.370 0.185 ;
        RECT  0.330 0.720 0.370 0.760 ;
        RECT  0.260 0.400 0.300 0.440 ;
        RECT  0.190 0.165 0.230 0.205 ;
        RECT  0.115 0.365 0.155 0.405 ;
        RECT  0.050 0.115 0.090 0.155 ;
        RECT  0.050 0.635 0.090 0.675 ;
        LAYER M1 ;
        RECT  0.405 0.380 0.435 0.460 ;
        RECT  0.355 0.240 0.405 0.655 ;
        RECT  0.250 0.240 0.355 0.290 ;
        RECT  0.095 0.605 0.355 0.655 ;
        RECT  0.170 0.145 0.250 0.290 ;
        RECT  0.045 0.605 0.095 0.695 ;
    END
END OR2SGD1BWP30P140




MACRO CKMUX2SGD1BWP30P140
    CLASS CORE ;
    FOREIGN CKMUX2SGD1BWP30P140 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 0.900 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.045475 ;
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  1.355 0.125 1.375 0.570 ;
        RECT  1.325 0.125 1.355 0.755 ;
        RECT  1.305 0.125 1.325 0.220 ;
        RECT  1.305 0.520 1.325 0.755 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.011100 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.345 0.155 0.445 ;
        RECT  0.045 0.345 0.115 0.555 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.010650 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M2 ;
        RECT  0.425 0.275 0.735 0.325 ;
        VIA  0.53 0.3 VIA12_square ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.011550 ;
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER M2 ;
        RECT  1.125 0.375 1.355 0.425 ;
        RECT  1.045 0.375 1.125 0.505 ;
        VIA  1.09 0.45 VIA12_square ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 -0.075 1.400 0.075 ;
        RECT  1.165 -0.075 1.215 0.180 ;
        RECT  0.510 -0.075 1.165 0.075 ;
        RECT  0.440 -0.075 0.510 0.195 ;
        RECT  0.095 -0.075 0.440 0.075 ;
        RECT  0.045 -0.075 0.095 0.180 ;
        RECT  0.000 -0.075 0.045 0.075 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 0.825 1.400 0.975 ;
        RECT  1.170 0.695 1.220 0.975 ;
        RECT  0.530 0.825 1.170 0.975 ;
        RECT  0.450 0.690 0.530 0.975 ;
        RECT  0.100 0.825 0.450 0.975 ;
        RECT  0.035 0.735 0.100 0.975 ;
        RECT  0.000 0.825 0.035 0.975 ;
        END
    END VDD
    OBS
        LAYER CO ;
        RECT  1.310 0.145 1.350 0.185 ;
        RECT  1.310 0.565 1.350 0.605 ;
        RECT  1.310 0.675 1.350 0.715 ;
        RECT  1.235 0.410 1.275 0.450 ;
        RECT  1.170 0.120 1.210 0.160 ;
        RECT  1.170 0.715 1.210 0.755 ;
        RECT  1.100 0.410 1.140 0.450 ;
        RECT  1.030 0.145 1.070 0.185 ;
        RECT  1.030 0.705 1.070 0.745 ;
        RECT  0.960 0.455 1.000 0.495 ;
        RECT  0.890 0.140 0.930 0.180 ;
        RECT  0.890 0.705 0.930 0.745 ;
        RECT  0.820 0.380 0.860 0.420 ;
        RECT  0.750 0.165 0.790 0.205 ;
        RECT  0.750 0.690 0.790 0.730 ;
        RECT  0.680 0.525 0.720 0.565 ;
        RECT  0.610 0.140 0.650 0.180 ;
        RECT  0.610 0.690 0.650 0.730 ;
        RECT  0.540 0.335 0.580 0.375 ;
        RECT  0.470 0.135 0.510 0.175 ;
        RECT  0.470 0.710 0.510 0.750 ;
        RECT  0.405 0.445 0.445 0.485 ;
        RECT  0.330 0.140 0.370 0.180 ;
        RECT  0.330 0.660 0.370 0.700 ;
        RECT  0.190 0.145 0.230 0.185 ;
        RECT  0.190 0.730 0.230 0.770 ;
        RECT  0.115 0.375 0.155 0.415 ;
        RECT  0.050 0.105 0.090 0.145 ;
        RECT  0.050 0.755 0.090 0.795 ;
        LAYER M1 ;
        RECT  1.255 0.390 1.275 0.470 ;
        RECT  1.205 0.275 1.255 0.625 ;
        RECT  0.800 0.275 1.205 0.325 ;
        RECT  0.930 0.575 1.205 0.625 ;
        RECT  1.055 0.375 1.155 0.525 ;
        RECT  0.980 0.675 1.120 0.775 ;
        RECT  1.000 0.135 1.115 0.225 ;
        RECT  0.955 0.435 1.005 0.525 ;
        RECT  0.870 0.135 1.000 0.185 ;
        RECT  0.810 0.475 0.955 0.525 ;
        RECT  0.860 0.575 0.930 0.765 ;
        RECT  0.710 0.375 0.880 0.425 ;
        RECT  0.760 0.475 0.810 0.575 ;
        RECT  0.595 0.675 0.805 0.745 ;
        RECT  0.750 0.145 0.800 0.325 ;
        RECT  0.710 0.525 0.760 0.575 ;
        RECT  0.660 0.375 0.710 0.475 ;
        RECT  0.660 0.525 0.710 0.625 ;
        RECT  0.560 0.125 0.700 0.225 ;
        RECT  0.515 0.425 0.660 0.475 ;
        RECT  0.385 0.575 0.660 0.625 ;
        RECT  0.455 0.275 0.600 0.375 ;
        RECT  0.405 0.425 0.515 0.525 ;
        RECT  0.355 0.125 0.385 0.195 ;
        RECT  0.355 0.575 0.385 0.720 ;
        RECT  0.305 0.125 0.355 0.720 ;
        RECT  0.205 0.125 0.255 0.775 ;
        RECT  0.170 0.125 0.205 0.225 ;
        RECT  0.170 0.725 0.205 0.775 ;
        LAYER VIA1 ;
        RECT  1.035 0.175 1.085 0.225 ;
        RECT  1.025 0.675 1.075 0.725 ;
        RECT  0.725 0.675 0.775 0.725 ;
        RECT  0.620 0.175 0.670 0.225 ;
        RECT  0.435 0.475 0.485 0.525 ;
        RECT  0.205 0.575 0.255 0.625 ;
        LAYER M2 ;
        RECT  0.985 0.175 1.115 0.225 ;
        RECT  0.985 0.675 1.105 0.725 ;
        RECT  0.935 0.175 0.985 0.725 ;
        RECT  0.835 0.175 0.885 0.725 ;
        RECT  0.590 0.175 0.835 0.225 ;
        RECT  0.695 0.675 0.835 0.725 ;
        RECT  0.425 0.445 0.495 0.625 ;
        RECT  0.155 0.575 0.425 0.625 ;
    END
END CKMUX2SGD1BWP30P140
